//TOP.v
module TOP(CLK, RST, EN);

input CLK, RST, EN;

//GOTO_ADDR.v
wire [11:0] ADDR_G;

//GOTO_RAM.v
wire [7:0] CURRENT_STATE_G, NEXT_STATE;//G=GOTO_FUNCTION
wire [3:0] CHARA;

//FAILURE_ADDR.v
wire [11:0] ADDR_F;

//FAILURE_RAM.v
wire [7:0] CURRENT_STATE_F, FAILURE_STATE;//F=FAILURE_FUNCITON

//TABLE_READER.v
wire [7:0] READER;
wire [7:0] READER1;
wire [7:0] RESULT;

GOTO_RAM GOTO_RAM(
    .CLK(CLK),
    .RST(RST), 
    .ADDR_G(ADDR_G),
    .CURRENT_STATE_G(CURRENT_STATE_G),
    .CHARA(CHARA),
    .NEXT_STATE(NEXT_STATE)
);

GOTO_ADDR GOTO_ADDR(
    .CLK(CLK),
    .RST(RST),
    .ADDR_G(ADDR_G)
);

FAILURE_RAM FAILURE_RAM(
    .CLK(CLK),
    .RST(RST), 
    .ADDR_F(ADDR_F),
    .CURRENT_STATE_F(CURRENT_STATE_F),
    .FAILURE_STATE(FAILURE_STATE)
);

FAILURE_ADDR FAILURE_ADDR(
    .CLK(CLK),
    .RST(RST),
    .ADDR_F(ADDR_F)
);

TABLE_READER TABLE_READER(
  .CLK(CLK),
  .RST(RST),
  .EN(EN),
  .READER(READER),
  .READER1(READER1),
  .RESULT(RESULT)
);

endmodule
